`include "uvm_macros.svh"

package fifo_pkg;
  import uvm_pkg::*;

  `include "defines_fifo.sv"

  `include "write_sequence_item_fifo.sv"
  `include "read_sequence_item_fifo.sv"

  `include "write_sequence_fifo.sv"
  `include "read_sequence_fifo.sv"

  `include "write_sequencer_fifo.sv"
  `include "read_sequencer_fifo.sv"

  `include "write_driver_fifo.sv"
  `include "read_driver_fifo.sv"

  `include "write_monitor_fifo.sv"
  `include "read_monitor_fifo.sv"

  `include "write_agent_fifo.sv"
  `include "read_agent_fifo.sv"

  `include "subscriber_fifo.sv"
  `include "scoreboard_fifo.sv"

  `include "virtual_sequencer_fifo.sv"
  `include "virtual_sequence_fifo.sv"

  `include "environment_fifo.sv"
  `include "test_fifo.sv"

endpackage

