
`define ADDR_WIDTH 4
`define DATA_WIDTH 8
`define no_of_trans 100
